module name();
initial begin
$display("My name is Hieu and I start the course today June 22th 2025");
end
endmodule

